library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package head_const is
	constant mul_delay: integer := 3;
	constant div_delay: integer := 4;
	constant fun_delay: integer := 2;
	constant fifo_delay: integer := 0;
end;

package body head_const is
end;
